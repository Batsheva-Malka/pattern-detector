// Pattern Detector Sequencer
// Standard UVM sequencer for pattern_detector_seq_item

typedef uvm_sequencer#(pattern_detector_seq_item) pattern_detector_sequencer;
